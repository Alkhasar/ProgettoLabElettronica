/**
*   Top Module for the CCD array DAQ
*
*   clk (wire in): Main FPGA clock
*   rst (wire in): Main async reset
*/

`timescale 10ns / 1ns

module Top (
    input wire clk,
    input wire rst
);

endmodule
